package axi_test_reg_rtl_pkg;
  localparam int REGISTER_0_BYTE_WIDTH = 4;
  localparam int REGISTER_0_BYTE_SIZE = 4;
  localparam bit [7:0] REGISTER_0_BYTE_OFFSET = 8'h00;
  localparam int REGISTER_0_BIT_FIELD_0_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_0_BIT_FIELD_0_BIT_MASK = 4'hf;
  localparam int REGISTER_0_BIT_FIELD_0_BIT_OFFSET = 0;
  localparam int REGISTER_0_BIT_FIELD_1_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_0_BIT_FIELD_1_BIT_MASK = 4'hf;
  localparam int REGISTER_0_BIT_FIELD_1_BIT_OFFSET = 4;
  localparam int REGISTER_0_BIT_FIELD_2_BIT_WIDTH = 1;
  localparam bit REGISTER_0_BIT_FIELD_2_BIT_MASK = 1'h1;
  localparam int REGISTER_0_BIT_FIELD_2_BIT_OFFSET = 8;
  localparam int REGISTER_0_BIT_FIELD_3_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_0_BIT_FIELD_3_BIT_MASK = 2'h3;
  localparam int REGISTER_0_BIT_FIELD_3_BIT_OFFSET = 9;
  localparam int REGISTER_0_BIT_FIELD_4_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_0_BIT_FIELD_4_BIT_MASK = 2'h3;
  localparam int REGISTER_0_BIT_FIELD_4_BIT_OFFSET = 11;
  localparam int REGISTER_0_BIT_FIELD_5_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_0_BIT_FIELD_5_BIT_MASK = 2'h3;
  localparam int REGISTER_0_BIT_FIELD_5_BIT_OFFSET = 13;
  localparam int REGISTER_0_BIT_FIELD_6_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_0_BIT_FIELD_6_BIT_MASK = 2'h3;
  localparam int REGISTER_0_BIT_FIELD_6_BIT_OFFSET = 15;
  localparam int REGISTER_1_BYTE_WIDTH = 4;
  localparam int REGISTER_1_BYTE_SIZE = 4;
  localparam bit [7:0] REGISTER_1_BYTE_OFFSET = 8'h04;
  localparam int REGISTER_1_BIT_WIDTH = 1;
  localparam bit REGISTER_1_BIT_MASK = 1'h1;
  localparam int REGISTER_1_BIT_OFFSET = 0;
  localparam bit REGISTER_1_FOO = 1'h0;
  localparam bit REGISTER_1_BAR = 1'h1;
  localparam int REGISTER_2_BYTE_WIDTH = 4;
  localparam int REGISTER_2_BYTE_SIZE = 4;
  localparam bit [7:0] REGISTER_2_BYTE_OFFSET = 8'h08;
  localparam int REGISTER_2_BIT_FIELD_0_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_2_BIT_FIELD_0_BIT_MASK = 4'hf;
  localparam int REGISTER_2_BIT_FIELD_0_BIT_OFFSET = 0;
  localparam int REGISTER_2_BIT_FIELD_1_BIT_WIDTH = 8;
  localparam bit [7:0] REGISTER_2_BIT_FIELD_1_BIT_MASK = 8'hff;
  localparam int REGISTER_2_BIT_FIELD_1_BIT_OFFSET = 8;
  localparam int REGISTER_2_BIT_FIELD_2_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_2_BIT_FIELD_2_BIT_MASK = 4'hf;
  localparam int REGISTER_2_BIT_FIELD_2_BIT_OFFSET = 16;
endpackage
